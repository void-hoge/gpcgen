module gpc1_1(input wire[0:0]src0, output wire[0:0]dst);
    assign dst[0] = src0[0];
endmodule

